module seg_secmin (
    input [5:0]value,
    output reg [6:0]seg0, seg1 // seg1: chuc, seg0: dv
);
    
    always @(value) begin
        case (value)

            0: {seg1, seg0} = 14'b0000001_0000001;
            1: {seg1, seg0} = 14'b0000001_1001111;
            2: {seg1, seg0} = 14'b0000001_0010010;
            3: {seg1, seg0} = 14'b0000001_0000110;
            4: {seg1, seg0} = 14'b0000001_1001100;
            5: {seg1, seg0} = 14'b0000001_0100100;
            6: {seg1, seg0} = 14'b0000001_0100000;
            7: {seg1, seg0} = 14'b0000001_0001111;
            8: {seg1, seg0} = 14'b0000001_0000000;
            9: {seg1, seg0} = 14'b0000001_0000100;

            10: {seg1, seg0} = 14'b1001111_0000001;
            11: {seg1, seg0} = 14'b1001111_1001111;
            12: {seg1, seg0} = 14'b1001111_0010010;
            13: {seg1, seg0} = 14'b1001111_0000110;
            14: {seg1, seg0} = 14'b1001111_1001100;
            15: {seg1, seg0} = 14'b1001111_0100100;
            16: {seg1, seg0} = 14'b1001111_0100000;
            17: {seg1, seg0} = 14'b1001111_0001111;
            18: {seg1, seg0} = 14'b1001111_0000000;
            19: {seg1, seg0} = 14'b1001111_0000100;

            20: {seg1, seg0} = 14'b0010010_0000001;
            21: {seg1, seg0} = 14'b0010010_1001111;
            22: {seg1, seg0} = 14'b0010010_0010010;
            23: {seg1, seg0} = 14'b0010010_0000110;
            24: {seg1, seg0} = 14'b0010010_1001100;
            25: {seg1, seg0} = 14'b0010010_0100100;
            26: {seg1, seg0} = 14'b0010010_0100000;
            27: {seg1, seg0} = 14'b0010010_0001111;
            28: {seg1, seg0} = 14'b0010010_0000000;
            29: {seg1, seg0} = 14'b0010010_0000100;

            30: {seg1, seg0} = 14'b0000110_0000001;
            31: {seg1, seg0} = 14'b0000110_1001111;
            32: {seg1, seg0} = 14'b0000110_0010010;
            33: {seg1, seg0} = 14'b0000110_0000110;
            34: {seg1, seg0} = 14'b0000110_1001100;
            35: {seg1, seg0} = 14'b0000110_0100100;
            36: {seg1, seg0} = 14'b0000110_0100000;
            37: {seg1, seg0} = 14'b0000110_0001111;
            38: {seg1, seg0} = 14'b0000110_0000000;
            39: {seg1, seg0} = 14'b0000110_0000100;

            40: {seg1, seg0} = 14'b1001100_0000001;
            41: {seg1, seg0} = 14'b1001100_1001111;
            42: {seg1, seg0} = 14'b1001100_0010010;
            43: {seg1, seg0} = 14'b1001100_0000110;
            44: {seg1, seg0} = 14'b1001100_1001100;
            45: {seg1, seg0} = 14'b1001100_0100100;
            46: {seg1, seg0} = 14'b1001100_0100000;
            47: {seg1, seg0} = 14'b1001100_0001111;
            48: {seg1, seg0} = 14'b1001100_0000000;
            49: {seg1, seg0} = 14'b1001100_0000100;

            50: {seg1, seg0} = 14'b0100100_0000001;
            51: {seg1, seg0} = 14'b0100100_1001111;
            52: {seg1, seg0} = 14'b0100100_0010010;
            53: {seg1, seg0} = 14'b0100100_0000110;
            54: {seg1, seg0} = 14'b0100100_1001100;
            55: {seg1, seg0} = 14'b0100100_0100100;
            56: {seg1, seg0} = 14'b0100100_0100000;
            57: {seg1, seg0} = 14'b0100100_0001111;
            58: {seg1, seg0} = 14'b0100100_0000000;
            59: {seg1, seg0} = 14'b0100100_0000100;

            default: {seg1, seg0} = 14'b1111111_1111111;
        endcase
    end

endmodule